`timescale 1ns / 1ps

`define ADD 4'b0000             
`define SUB 4'b1000             
`define SLL 4'b0001             
`define SRL 4'b0101             
`define SRA 4'b1101 
`define SLT 4'b0010 
`define SLU 4'b0011
`define XOR 4'b0100
`define OR  4'b0110
`define AND 4'b0111

`define OP_TYPE_R 7'b0110011