`timescale 1ns / 1ps
`include "defines.sv"

module ControlUnit (
    input  logic [31:0] instrCode,
    output logic        regFileWe,
    output logic        aluSrcMuxSel,
    output logic [ 3:0] aluControl,
    output logic        busWe,
    output logic [ 2:0] RFWDSrcMuxSel,
    output logic        branch,
    output logic        JAL,
    output logic        JALR
);
    wire  [6:0] opcode = instrCode[6:0];
    wire  [3:0] operator = {instrCode[30], instrCode[14:12]};
    logic [8:0] signals;

    assign {regFileWe, aluSrcMuxSel, busWe, RFWDSrcMuxSel, branch, JAL, JALR} = signals;

    always_comb begin
        signals = 0;
        case (opcode)
            //{regFileWe, aluSrcMuxSel, busWe, RFWDSrcMuxSel, branch, JAL, JALR}
            `OP_TYPE_R:     signals = 9'b1_0_0_000_0_0_0;
            `OP_TYPE_I:     signals = 9'b1_1_0_000_0_0_0;
            `OP_TYPE_S:     signals = 9'b0_1_1_000_0_0_0;
            `OP_TYPE_L:     signals = 9'b1_1_0_001_0_0_0;
            `OP_TYPE_B:     signals = 9'b0_0_0_000_1_0_0;
            `OP_TYPE_JAL:   signals = 9'b1_0_0_010_0_1_0;
            `OP_TYPE_JALR:  signals = 9'b1_0_0_010_0_0_1;
            `OP_TYPE_LUI:   signals = 9'b1_0_0_011_0_0_0;
            `OP_TYPE_AUIPC: signals = 9'b1_0_0_100_0_0_0;
            default:        signals = 0;
        endcase
    end

    always_comb begin
        aluControl = `ADD;
        case (opcode)
            `OP_TYPE_R:    aluControl = operator;
            `OP_TYPE_B:    aluControl = operator;
            `OP_TYPE_JAL:  aluControl = operator;
            `OP_TYPE_JALR: aluControl = operator;
            //`OP_TYPE_S: aluControl = operator; default 출력으로 나가도록 함.
            `OP_TYPE_I: begin
                if (operator == 4'b1101) aluControl = operator;
                else aluControl = {1'b0, operator[2:0]};
            end
            default:       aluControl = `ADD;
        endcase
    end

endmodule
